module top(
   input logic btnu, student, prof, pm,
   input logic[3:0] hour,
   input logic[8:0] sw,
   output logic[15:0] led
);

//Code Goes Here

endmodule
