module top(
   input logic[15:0] sw,
   input logic btnl,
   output logic[15:0] led
);

//Code Goes Here

endmodule
