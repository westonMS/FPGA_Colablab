module add_8(
  input logic Cin,
  input logic [7:0] a, b,
  output logic [7:0] s,
  output logic Cout 
  );
  //Instantiate 8 instances of full_adder
  //Have Cin be the first carry in and Cout be the last carry out
  
 endmodule
