module full_add(
  input logic a, b, Cin,
  output logic s, Cout
  );
  //A, B and the Cin should be added together. s is the result and Cout signifies carry over.
  endmodule
