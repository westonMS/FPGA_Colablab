module top(
   input logic[12:0] sw,
   input logic btnr, A, B, C,
   output logic[15:0] led
);

//Code Goes Here

endmodule
